`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Extend the data (2->8)
//////////////////////////////////////////////////////////////////////////////////
module sign_extender(
    input [1:0] in,
    output [7:0] out
    );
	 
	assign out = (in[1] ? {6'b111111, in[1:0]} : {6'b000000, in[1:0]});
	
endmodule